// Control Block
module control(
    input [5:0] opcode,
    output regDest,
    output jump,
    output branch,
    output memRead,
    output memToReg,
    output aluOp,
    output memWrite,
    output aluSrc,
    output regWrite
);




endmodule